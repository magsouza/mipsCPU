module MUX3 (WriteData, w_ALUResult, w_SS, w_MUX3);

	input WriteData;
	input [31:0] w_ALUResult, w_SS;
	output reg[31:0] w_MUX3;

always @(*)

begin
	case (WriteData)
		1'b0: begin
			w_MUX3[31:0] <= w_ALUResult[31:0];
		end
		1'b1: begin
			w_MUX3[31:0] <= w_SS[31:0];
		end
	endcase
end

endmodule
